module chessController(input  logic signal,
                       output logic)
