/*
Encoding:
color: black = 1, white = 0
position (0,0) is in top left of board
position (7,7) is in bottom right of board
rook allowable moves: 
rookAllowUp[2:0]
rookAllowRight[2:0]
rookAllowDown[2:0]
rookAllowLeft[2:0]
*/
